netcdf weak_monotonic_coordinate {

dimensions:
    lon = 3 ;
    lat = 3 ;
    time1 = 3 ;
    time2 = 3 ;
    time3 = 3 ;

variables:
    // weak-monotonic coordinate.
    int wind1(time1, lat, lon) ;
        wind1:standard_name = "eastward_wind" ;
        wind1:units = "m s-1" ;
        wind1:test = "weak-monotonic time coordinate" ;

    // masked monotonic coordinate.
    int wind2(time2, lat, lon) ;
        wind2:standard_name = "eastward_wind" ;
        wind2:units = "m s-1" ;
        wind2:test = "masked monotonic time coordinate" ;

    // masked non-monotonic coordinate.
    int wind3(time3, lat, lon) ;
        wind3:standard_name = "eastward_wind" ;
        wind3:units = "m s-1" ;
        wind3:test = "masked non-monotonic time coordinate" ;

    int lon(lon) ;
        lon:standard_name = "longitude" ;
        lon:units = "degrees_east" ;

    int lat(lat) ;
        lat:standard_name = "latitude" ;
        lat:units = "degrees_north" ;

    // weak-monotonic coordinate.
    int time1(time1) ;
        time1:standard_name = "time" ;
        time1:units = "hours since 1970-01-01 00:00:00" ;

    // masked monotonic coordinate.
    int time2(time2) ;
        time2:standard_name = "time" ;
        time2:units = "hours since 1970-01-01 00:00:00" ;
        time2:_FillValue = 100 ;
 
    // masked non-monotonic coordinate.
    int time3(time3) ;
        time3:standard_name = "time" ;
        time3:units = "hours since 1970-01-01 00:00:00" ;   
        time3:_FillValue = 100 ;

data:
    wind1 = 1,  2,  3,  4,  5,  6,  7,  8,  9,
            10, 11, 12, 13, 14, 15, 16, 17, 18,
            19, 20, 21, 22, 23, 24, 25, 26, 27 ;

    wind2 = 1,  2,  3,  4,  5,  6,  7,  8,  9,
            10, 11, 12, 13, 14, 15, 16, 17, 18,
            19, 20, 21, 22, 23, 24, 25, 26, 27 ;

    wind2 = 1,  2,  3,  4,  5,  6,  7,  8,  9,
            10, 11, 12, 13, 14, 15, 16, 17, 18,
            19, 20, 21, 22, 23, 24, 25, 26, 27 ;

    lon = 10, 20, 30, 40, 50 ;

    lat = 50, 60, 70, 80 ;

    // weak-monotonic coordinate.
    time1 = 1, 1, 2 ;

    // masked monotonic coordinate.
    time2 = 1, 2, _ ;

    // masked non-monotonic coordinate.
    time3 = 1, _, 3 ;

}
